-------------------------------------------------------------------------------
--
-- ✄╔╗──╔╗╔╗───╔╗╔╗
-- ✄║║──║║║║───║║║║
-- ✄║║╔╦╣║║║╔══╣║║║─╔╦══╗
-- ✄║╚╝╬╣║║║║╔╗║║║║─╠╣╔╗║
-- ✄║╔╗╣║╚╣╚╣╔╗║╚╣╚╦╣║╚╝║
-- ✄╚╝╚╩╩═╩═╩╝╚╩═╩═╩╩╩══╝
--
-------------------------------------------------------------------------------
--
-- Company: killall.io
-- Author: Joachim Schmidt <joachim.schmidt@semaphore-networks.ch
--
-- Module Name: tb_killallio_sig_sync - arch
-- Target Device: hepia-cores.ch:scalp_node:part0:0.1 xc7z015clg485-2
-- Tool version: 2022.1
-- Description: Testbench for killallio_sig_sync
--
-- Last update: 2022-06-08
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_killallio_sig_sync is
end tb_killallio_sig_sync;

architecture behavioral of tb_killallio_sig_sync is

begin

end behavioral;
